// mcp program to debug UART 

  $display("UART_DEBUG.MCP RUNNING");
