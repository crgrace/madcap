///////////////////////////////////////////////////////////////////
// File Name: gate_posedge_clk.sv
// Engineer:  Dario Gnani (dgnani@lbl.gov)
// Description: Clock gating logic for posedge-sensitive seq logic.
//              Basic description of integrated clock gating (ICG) cell.
//
// NOTE: pin names must be EN, TE, CLK, ENCLK (!)
///////////////////////////////////////////////////////////////////
`timescale 1ns / 10ps
module gate_posedge_clk
    (output logic ENCLK,           // gated posedge clock
    input logic EN,               // clock-gating: enable clock (active high)
    input logic CLK);             // posedge clock

/* //DG: could not map correctly!? 
// Internal Variables 
logic Esync;

// UART TX Logic
always_latch  
    if (!CLK)
        Esync <= EN; 
    // always_latch

always_comb
   ENCLK = Esync & CLK;
*/
/*//DG: could not map correctly!?
always_latch  
    if (!CLK)
	if (EN)
           ENCLK <= CLK; 
    // always_latch
*/
logic EN_dly;
always @(EN) EN_dly = #1.5 EN; //DG: required to suppress timing violations
//this is clearly acceptable only if the EN is generated by the same clock we are gating

//TP: updated to 130nm gated clock latch
/*TLATNCAX8 
    mapped_ICGP(
    .ECK(ENCLK),
    .E(EN_dly),
    .CK(CLK)
    );
*/
CKLNQD8
    mapped_ICGP(
    .Q(ENCLK),
    .TE(1'b0),
    .E(EN_dly),
    .CP(CLK)
    );

endmodule

